module i2c_phy_bit_ctl(
    input   clk,
    input   rstn,

    input   [2:0]   cmd,
    output          ack,
    input           scl_i,
    input           sda_i,
    output          scl_o,
    output          sda_o
);






endmodule
