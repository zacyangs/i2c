interface interrupt(input clk);

    logic irq_gold;
    logic irq_dut;

endinterface
