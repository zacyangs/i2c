package pkg;
    `include "./test_case/test_base.sv"
    `include "./test_case/test_reg.sv"
    `include "./test_case/test_slv.sv"
    `include "factory.sv"
    `include "env.sv"
endpackage
